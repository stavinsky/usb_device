module queue #(parameter size = 256) (r_clk, data_out, w_clk, data_in, empty, full, rst, r_en, w_en);
    input wire r_clk;
    output [7:0]data_out;

    input wire w_clk;
    input [7:0]data_in;

    output empty;
    output full;
    input rst;
    input r_en;
    input w_en;

    localparam adr_size = $clog2(size) -1 ;
    (* ram_style = "block" *)
    reg [7:0] mem [0:size-1];
    reg [adr_size:0] r_address = 0;
    reg [adr_size:0] w_address = 0;

    // assign data_out = mem[r_address];
    reg [7:0] r_data_out;
    assign data_out = r_data_out;
    always @(posedge r_clk or negedge rst) begin
        if (~rst) begin
            r_address <= 0;
        end
        else if (~empty && r_en) begin
            r_address <= r_address + 1'b1;
        end
    end
    wire clk;
    assign clk = r_clk | w_clk;
    always @(posedge clk) begin
         r_data_out <= mem[r_address];
    end
    always @(posedge w_clk or negedge rst) begin
        if (~rst) begin
            w_address <= 0;
        end
        else if  (~full && w_en) begin
            w_address <= w_address + 1'b1;
        end
    end
    always @(posedge w_clk ) begin
        if  (~full && w_en) begin
            mem[w_address] <= data_in;
        end
    end
    assign empty = r_address == w_address;
    assign full = (w_address + 1'b1) == r_address;
endmodule
